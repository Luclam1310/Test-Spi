package spi_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "tb_defines.svh"
`include "spi_seq_item.svh"
`include "wb_bfm.svh"
`include "spi_driver.svh"
`include "spi_monitor.svh"
`include "spi_sequencer.svh"
`include "spi_agent.svh"
`include "spi_coverage.svh"
`include "spi_scoreboard.svh"
`include "spi_seq.svh"
`include "spi_env.svh"
`include "spi_test.svh"

endpackage 

